LIBRARY IEEE;
USE ieee.std_logic_1164.ALL;

PACKAGE array_integer IS
	--GENERIC( data_width : INTEGER := 10);
	TYPE integer_array IS ARRAY(9 DOWNTO 0) OF integer;

END array_integer;

PACKAGE BODY array_integer IS
END array_integer;