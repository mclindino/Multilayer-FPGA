LIBRARY IEEE;
USE ieee.std_logic_1164.ALL;
USE work.parameters.ALL;

ENTITY max_pooling IS
PORT(
		input		: IN  array_neuron;
		output	: OUT array_neuron
);
END max_pooling;

ARCHITECTURE behavior OF max_pooling IS
BEGIN

END behavior;